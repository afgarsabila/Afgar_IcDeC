magic
tech sky130A
magscale 1 2
timestamp 1729133440
<< nwell >>
rect -296 -1373 296 1373
<< pmos >>
rect -100 754 100 1154
rect -100 118 100 518
rect -100 -518 100 -118
rect -100 -1154 100 -754
<< pdiff >>
rect -158 1142 -100 1154
rect -158 766 -146 1142
rect -112 766 -100 1142
rect -158 754 -100 766
rect 100 1142 158 1154
rect 100 766 112 1142
rect 146 766 158 1142
rect 100 754 158 766
rect -158 506 -100 518
rect -158 130 -146 506
rect -112 130 -100 506
rect -158 118 -100 130
rect 100 506 158 518
rect 100 130 112 506
rect 146 130 158 506
rect 100 118 158 130
rect -158 -130 -100 -118
rect -158 -506 -146 -130
rect -112 -506 -100 -130
rect -158 -518 -100 -506
rect 100 -130 158 -118
rect 100 -506 112 -130
rect 146 -506 158 -130
rect 100 -518 158 -506
rect -158 -766 -100 -754
rect -158 -1142 -146 -766
rect -112 -1142 -100 -766
rect -158 -1154 -100 -1142
rect 100 -766 158 -754
rect 100 -1142 112 -766
rect 146 -1142 158 -766
rect 100 -1154 158 -1142
<< pdiffc >>
rect -146 766 -112 1142
rect 112 766 146 1142
rect -146 130 -112 506
rect 112 130 146 506
rect -146 -506 -112 -130
rect 112 -506 146 -130
rect -146 -1142 -112 -766
rect 112 -1142 146 -766
<< nsubdiff >>
rect -260 1303 -164 1337
rect 164 1303 260 1337
rect -260 1241 -226 1303
rect 226 1241 260 1303
rect -260 -1303 -226 -1241
rect 226 -1303 260 -1241
rect -260 -1337 -164 -1303
rect 164 -1337 260 -1303
<< nsubdiffcont >>
rect -164 1303 164 1337
rect -260 -1241 -226 1241
rect 226 -1241 260 1241
rect -164 -1337 164 -1303
<< poly >>
rect -100 1235 100 1251
rect -100 1201 -84 1235
rect 84 1201 100 1235
rect -100 1154 100 1201
rect -100 707 100 754
rect -100 673 -84 707
rect 84 673 100 707
rect -100 657 100 673
rect -100 599 100 615
rect -100 565 -84 599
rect 84 565 100 599
rect -100 518 100 565
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -118 100 -71
rect -100 -565 100 -518
rect -100 -599 -84 -565
rect 84 -599 100 -565
rect -100 -615 100 -599
rect -100 -673 100 -657
rect -100 -707 -84 -673
rect 84 -707 100 -673
rect -100 -754 100 -707
rect -100 -1201 100 -1154
rect -100 -1235 -84 -1201
rect 84 -1235 100 -1201
rect -100 -1251 100 -1235
<< polycont >>
rect -84 1201 84 1235
rect -84 673 84 707
rect -84 565 84 599
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -599 84 -565
rect -84 -707 84 -673
rect -84 -1235 84 -1201
<< locali >>
rect -260 1303 -164 1337
rect 164 1303 260 1337
rect -260 1241 -226 1303
rect 226 1241 260 1303
rect -100 1201 -84 1235
rect 84 1201 100 1235
rect -146 1142 -112 1158
rect -146 750 -112 766
rect 112 1142 146 1158
rect 112 750 146 766
rect -100 673 -84 707
rect 84 673 100 707
rect -100 565 -84 599
rect 84 565 100 599
rect -146 506 -112 522
rect -146 114 -112 130
rect 112 506 146 522
rect 112 114 146 130
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -130 -112 -114
rect -146 -522 -112 -506
rect 112 -130 146 -114
rect 112 -522 146 -506
rect -100 -599 -84 -565
rect 84 -599 100 -565
rect -100 -707 -84 -673
rect 84 -707 100 -673
rect -146 -766 -112 -750
rect -146 -1158 -112 -1142
rect 112 -766 146 -750
rect 112 -1158 146 -1142
rect -100 -1235 -84 -1201
rect 84 -1235 100 -1201
rect -260 -1303 -226 -1241
rect 226 -1303 260 -1241
rect -260 -1337 -164 -1303
rect 164 -1337 260 -1303
<< viali >>
rect -84 1201 84 1235
rect -146 766 -112 1142
rect 112 766 146 1142
rect -84 673 84 707
rect -84 565 84 599
rect -146 130 -112 506
rect 112 130 146 506
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -506 -112 -130
rect 112 -506 146 -130
rect -84 -599 84 -565
rect -84 -707 84 -673
rect -146 -1142 -112 -766
rect 112 -1142 146 -766
rect -84 -1235 84 -1201
<< metal1 >>
rect -96 1235 96 1241
rect -96 1201 -84 1235
rect 84 1201 96 1235
rect -96 1195 96 1201
rect -152 1142 -106 1154
rect -152 766 -146 1142
rect -112 766 -106 1142
rect -152 754 -106 766
rect 106 1142 152 1154
rect 106 766 112 1142
rect 146 766 152 1142
rect 106 754 152 766
rect -96 707 96 713
rect -96 673 -84 707
rect 84 673 96 707
rect -96 667 96 673
rect -96 599 96 605
rect -96 565 -84 599
rect 84 565 96 599
rect -96 559 96 565
rect -152 506 -106 518
rect -152 130 -146 506
rect -112 130 -106 506
rect -152 118 -106 130
rect 106 506 152 518
rect 106 130 112 506
rect 146 130 152 506
rect 106 118 152 130
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -130 -106 -118
rect -152 -506 -146 -130
rect -112 -506 -106 -130
rect -152 -518 -106 -506
rect 106 -130 152 -118
rect 106 -506 112 -130
rect 146 -506 152 -130
rect 106 -518 152 -506
rect -96 -565 96 -559
rect -96 -599 -84 -565
rect 84 -599 96 -565
rect -96 -605 96 -599
rect -96 -673 96 -667
rect -96 -707 -84 -673
rect 84 -707 96 -673
rect -96 -713 96 -707
rect -152 -766 -106 -754
rect -152 -1142 -146 -766
rect -112 -1142 -106 -766
rect -152 -1154 -106 -1142
rect 106 -766 152 -754
rect 106 -1142 112 -766
rect 146 -1142 152 -766
rect 106 -1154 152 -1142
rect -96 -1201 96 -1195
rect -96 -1235 -84 -1201
rect 84 -1235 96 -1201
rect -96 -1241 96 -1235
<< properties >>
string FIXED_BBOX -243 -1320 243 1320
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 1 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
