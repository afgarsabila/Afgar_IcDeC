magic
tech sky130A
magscale 1 2
timestamp 1729346457
<< nmos >>
rect -407 -131 -247 69
rect -189 -131 -29 69
rect 29 -131 189 69
rect 247 -131 407 69
<< ndiff >>
rect -465 57 -407 69
rect -465 -119 -453 57
rect -419 -119 -407 57
rect -465 -131 -407 -119
rect -247 57 -189 69
rect -247 -119 -235 57
rect -201 -119 -189 57
rect -247 -131 -189 -119
rect -29 57 29 69
rect -29 -119 -17 57
rect 17 -119 29 57
rect -29 -131 29 -119
rect 189 57 247 69
rect 189 -119 201 57
rect 235 -119 247 57
rect 189 -131 247 -119
rect 407 57 465 69
rect 407 -119 419 57
rect 453 -119 465 57
rect 407 -131 465 -119
<< ndiffc >>
rect -453 -119 -419 57
rect -235 -119 -201 57
rect -17 -119 17 57
rect 201 -119 235 57
rect 419 -119 453 57
<< poly >>
rect -407 141 -247 157
rect -407 107 -391 141
rect -263 107 -247 141
rect -407 69 -247 107
rect -189 141 -29 157
rect -189 107 -173 141
rect -45 107 -29 141
rect -189 69 -29 107
rect 29 141 189 157
rect 29 107 45 141
rect 173 107 189 141
rect 29 69 189 107
rect 247 141 407 157
rect 247 107 263 141
rect 391 107 407 141
rect 247 69 407 107
rect -407 -157 -247 -131
rect -189 -157 -29 -131
rect 29 -157 189 -131
rect 247 -157 407 -131
<< polycont >>
rect -391 107 -263 141
rect -173 107 -45 141
rect 45 107 173 141
rect 263 107 391 141
<< locali >>
rect -407 107 -391 141
rect -263 107 -247 141
rect -189 107 -173 141
rect -45 107 -29 141
rect 29 107 45 141
rect 173 107 189 141
rect 247 107 263 141
rect 391 107 407 141
rect -453 57 -419 73
rect -453 -135 -419 -119
rect -235 57 -201 73
rect -235 -135 -201 -119
rect -17 57 17 73
rect -17 -135 17 -119
rect 201 57 235 73
rect 201 -135 235 -119
rect 419 57 453 73
rect 419 -135 453 -119
<< viali >>
rect -391 107 -263 141
rect -173 107 -45 141
rect 45 107 173 141
rect 263 107 391 141
rect -453 -119 -419 57
rect -235 -119 -201 57
rect -17 -119 17 57
rect 201 -119 235 57
rect 419 -119 453 57
<< metal1 >>
rect -403 141 -251 147
rect -403 107 -391 141
rect -263 107 -251 141
rect -403 101 -251 107
rect -185 141 -33 147
rect -185 107 -173 141
rect -45 107 -33 141
rect -185 101 -33 107
rect 33 141 185 147
rect 33 107 45 141
rect 173 107 185 141
rect 33 101 185 107
rect 251 141 403 147
rect 251 107 263 141
rect 391 107 403 141
rect 251 101 403 107
rect -459 57 -413 69
rect -459 -119 -453 57
rect -419 -119 -413 57
rect -459 -131 -413 -119
rect -241 57 -195 69
rect -241 -119 -235 57
rect -201 -119 -195 57
rect -241 -131 -195 -119
rect -23 57 23 69
rect -23 -119 -17 57
rect 17 -119 23 57
rect -23 -131 23 -119
rect 195 57 241 69
rect 195 -119 201 57
rect 235 -119 241 57
rect 195 -131 241 -119
rect 413 57 459 69
rect 413 -119 419 57
rect 453 -119 459 57
rect 413 -131 459 -119
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.8 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
