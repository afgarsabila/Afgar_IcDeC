magic
tech sky130A
magscale 1 2
timestamp 1729362917
<< metal1 >>
rect -4692 2812 -537 2846
rect -4692 -1033 -4658 2812
rect -4397 2545 -1522 2602
rect -4397 1114 -4362 2545
rect -4071 2252 -4065 2304
rect -4013 2252 -4007 2304
rect -4056 1792 -4022 2252
rect -1555 2163 -1522 2545
rect -3881 2038 -2540 2082
rect -3881 1780 -3842 2038
rect -2574 1691 -2540 2038
rect -2115 1861 -2081 1908
rect -1555 1692 -1521 2163
rect -1113 1816 -1061 1822
rect -1113 1758 -1061 1764
rect -4398 1079 -4061 1114
rect -1983 290 -1939 415
rect -1985 210 -1939 290
rect -1985 95 -1941 210
rect -2903 51 -1941 95
rect -4055 -1033 -4021 -942
rect -4692 -1067 -4021 -1033
rect -2903 -1133 -2859 51
rect -1104 -206 -1070 1758
rect -571 1619 -537 2812
rect 582 2597 634 2603
rect 582 2539 634 2545
rect 72 1816 124 1822
rect 124 1773 324 1807
rect 72 1758 124 1764
rect 289 982 323 1773
rect 151 981 323 982
rect -129 948 323 981
rect -129 947 204 948
rect -283 770 321 804
rect -514 394 -446 476
rect -514 360 326 394
rect -514 359 -446 360
rect -1578 -240 -1070 -206
rect -1582 -868 -1034 -835
rect -1930 -1133 -1886 -966
rect -2903 -1177 -1886 -1133
rect -1067 -1162 -1034 -868
rect 591 -1162 624 2539
rect -1067 -1195 624 -1162
<< via1 >>
rect -4065 2252 -4013 2304
rect -1113 1764 -1061 1816
rect 582 2545 634 2597
rect 72 1764 124 1816
<< metal2 >>
rect -179 2542 -170 2602
rect -110 2588 -101 2602
rect 576 2588 582 2597
rect -110 2555 582 2588
rect -110 2542 -101 2555
rect 576 2545 582 2555
rect 634 2545 640 2597
rect -4065 2304 -4013 2310
rect -433 2308 -373 2317
rect -4013 2261 -433 2295
rect -4065 2246 -4013 2252
rect -433 2239 -373 2248
rect -1984 1764 -1937 2134
rect -1119 1764 -1113 1816
rect -1061 1807 -1055 1816
rect 66 1807 72 1816
rect -1061 1773 72 1807
rect -1061 1764 -1055 1773
rect 66 1764 72 1773
rect 124 1764 130 1816
rect -1984 1741 -1936 1764
rect -1983 1628 -1936 1741
<< via2 >>
rect -170 2542 -110 2602
rect -433 2248 -373 2308
<< metal3 >>
rect -175 2602 -105 2607
rect -175 2542 -170 2602
rect -110 2542 -105 2602
rect -175 2537 -105 2542
rect -438 2308 -366 2324
rect -438 2248 -433 2308
rect -373 2248 -366 2308
rect -438 1218 -366 2248
rect -171 1496 -109 2537
rect -437 1213 -373 1218
use nmos2  nmos2_0
timestamp 1729346615
transform 1 0 -2593 0 1 -571
box -208 -442 1155 528
use nmoscs  nmoscs_0
timestamp 1729234872
transform 1 0 -2387 0 1 1166
box -419 -772 1211 742
use pmos2  pmos2_0
timestamp 1729339022
transform 1 0 -622 0 1 930
box -335 -1922 810 746
use pmoscs  pmoscs_1
timestamp 1729355461
transform 1 0 -4015 0 1 -171
box -249 -833 916 2158
<< labels >>
flabel metal1 282 784 283 790 0 FreeSans 800 0 0 0 VIP
port 0 nsew
flabel metal1 259 378 259 378 0 FreeSans 800 0 0 0 VIN
port 1 nsew
flabel metal2 -1959 2098 -1959 2098 0 FreeSans 800 0 0 0 RS
port 2 nsew
flabel metal1 -550 1950 -550 1950 0 FreeSans 800 0 0 0 VDD
port 3 nsew
flabel metal1 -1961 257 -1961 257 0 FreeSans 800 0 0 0 GND
port 4 nsew
flabel metal3 -144 2424 -144 2424 0 FreeSans 800 0 0 0 OUT
port 5 nsew
<< end >>
