magic
tech sky130A
magscale 1 2
timestamp 1729133440
<< nwell >>
rect -396 -973 396 973
<< pmos >>
rect -200 554 200 754
rect -200 118 200 318
rect -200 -318 200 -118
rect -200 -754 200 -554
<< pdiff >>
rect -258 742 -200 754
rect -258 566 -246 742
rect -212 566 -200 742
rect -258 554 -200 566
rect 200 742 258 754
rect 200 566 212 742
rect 246 566 258 742
rect 200 554 258 566
rect -258 306 -200 318
rect -258 130 -246 306
rect -212 130 -200 306
rect -258 118 -200 130
rect 200 306 258 318
rect 200 130 212 306
rect 246 130 258 306
rect 200 118 258 130
rect -258 -130 -200 -118
rect -258 -306 -246 -130
rect -212 -306 -200 -130
rect -258 -318 -200 -306
rect 200 -130 258 -118
rect 200 -306 212 -130
rect 246 -306 258 -130
rect 200 -318 258 -306
rect -258 -566 -200 -554
rect -258 -742 -246 -566
rect -212 -742 -200 -566
rect -258 -754 -200 -742
rect 200 -566 258 -554
rect 200 -742 212 -566
rect 246 -742 258 -566
rect 200 -754 258 -742
<< pdiffc >>
rect -246 566 -212 742
rect 212 566 246 742
rect -246 130 -212 306
rect 212 130 246 306
rect -246 -306 -212 -130
rect 212 -306 246 -130
rect -246 -742 -212 -566
rect 212 -742 246 -566
<< nsubdiff >>
rect -360 903 -264 937
rect 264 903 360 937
rect -360 841 -326 903
rect 326 841 360 903
rect -360 -903 -326 -841
rect 326 -903 360 -841
rect -360 -937 -264 -903
rect 264 -937 360 -903
<< nsubdiffcont >>
rect -264 903 264 937
rect -360 -841 -326 841
rect 326 -841 360 841
rect -264 -937 264 -903
<< poly >>
rect -200 835 200 851
rect -200 801 -184 835
rect 184 801 200 835
rect -200 754 200 801
rect -200 507 200 554
rect -200 473 -184 507
rect 184 473 200 507
rect -200 457 200 473
rect -200 399 200 415
rect -200 365 -184 399
rect 184 365 200 399
rect -200 318 200 365
rect -200 71 200 118
rect -200 37 -184 71
rect 184 37 200 71
rect -200 21 200 37
rect -200 -37 200 -21
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -200 -118 200 -71
rect -200 -365 200 -318
rect -200 -399 -184 -365
rect 184 -399 200 -365
rect -200 -415 200 -399
rect -200 -473 200 -457
rect -200 -507 -184 -473
rect 184 -507 200 -473
rect -200 -554 200 -507
rect -200 -801 200 -754
rect -200 -835 -184 -801
rect 184 -835 200 -801
rect -200 -851 200 -835
<< polycont >>
rect -184 801 184 835
rect -184 473 184 507
rect -184 365 184 399
rect -184 37 184 71
rect -184 -71 184 -37
rect -184 -399 184 -365
rect -184 -507 184 -473
rect -184 -835 184 -801
<< locali >>
rect -360 903 -264 937
rect 264 903 360 937
rect -360 841 -326 903
rect 326 841 360 903
rect -200 801 -184 835
rect 184 801 200 835
rect -246 742 -212 758
rect -246 550 -212 566
rect 212 742 246 758
rect 212 550 246 566
rect -200 473 -184 507
rect 184 473 200 507
rect -200 365 -184 399
rect 184 365 200 399
rect -246 306 -212 322
rect -246 114 -212 130
rect 212 306 246 322
rect 212 114 246 130
rect -200 37 -184 71
rect 184 37 200 71
rect -200 -71 -184 -37
rect 184 -71 200 -37
rect -246 -130 -212 -114
rect -246 -322 -212 -306
rect 212 -130 246 -114
rect 212 -322 246 -306
rect -200 -399 -184 -365
rect 184 -399 200 -365
rect -200 -507 -184 -473
rect 184 -507 200 -473
rect -246 -566 -212 -550
rect -246 -758 -212 -742
rect 212 -566 246 -550
rect 212 -758 246 -742
rect -200 -835 -184 -801
rect 184 -835 200 -801
rect -360 -903 -326 -841
rect 326 -903 360 -841
rect -360 -937 -264 -903
rect 264 -937 360 -903
<< viali >>
rect -184 801 184 835
rect -246 566 -212 742
rect 212 566 246 742
rect -184 473 184 507
rect -184 365 184 399
rect -246 130 -212 306
rect 212 130 246 306
rect -184 37 184 71
rect -184 -71 184 -37
rect -246 -306 -212 -130
rect 212 -306 246 -130
rect -184 -399 184 -365
rect -184 -507 184 -473
rect -246 -742 -212 -566
rect 212 -742 246 -566
rect -184 -835 184 -801
<< metal1 >>
rect -196 835 196 841
rect -196 801 -184 835
rect 184 801 196 835
rect -196 795 196 801
rect -252 742 -206 754
rect -252 566 -246 742
rect -212 566 -206 742
rect -252 554 -206 566
rect 206 742 252 754
rect 206 566 212 742
rect 246 566 252 742
rect 206 554 252 566
rect -196 507 196 513
rect -196 473 -184 507
rect 184 473 196 507
rect -196 467 196 473
rect -196 399 196 405
rect -196 365 -184 399
rect 184 365 196 399
rect -196 359 196 365
rect -252 306 -206 318
rect -252 130 -246 306
rect -212 130 -206 306
rect -252 118 -206 130
rect 206 306 252 318
rect 206 130 212 306
rect 246 130 252 306
rect 206 118 252 130
rect -196 71 196 77
rect -196 37 -184 71
rect 184 37 196 71
rect -196 31 196 37
rect -196 -37 196 -31
rect -196 -71 -184 -37
rect 184 -71 196 -37
rect -196 -77 196 -71
rect -252 -130 -206 -118
rect -252 -306 -246 -130
rect -212 -306 -206 -130
rect -252 -318 -206 -306
rect 206 -130 252 -118
rect 206 -306 212 -130
rect 246 -306 252 -130
rect 206 -318 252 -306
rect -196 -365 196 -359
rect -196 -399 -184 -365
rect 184 -399 196 -365
rect -196 -405 196 -399
rect -196 -473 196 -467
rect -196 -507 -184 -473
rect 184 -507 196 -473
rect -196 -513 196 -507
rect -252 -566 -206 -554
rect -252 -742 -246 -566
rect -212 -742 -206 -566
rect -252 -754 -206 -742
rect 206 -566 252 -554
rect 206 -742 212 -566
rect 246 -742 252 -566
rect 206 -754 252 -742
rect -196 -801 196 -795
rect -196 -835 -184 -801
rect 184 -835 196 -801
rect -196 -841 196 -835
<< properties >>
string FIXED_BBOX -343 -920 343 920
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 2 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
