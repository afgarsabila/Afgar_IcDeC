magic
tech sky130A
magscale 1 2
timestamp 1729234872
<< psubdiff >>
rect -419 695 -359 729
rect 1151 695 1211 729
rect -419 669 -385 695
rect 1177 669 1211 695
rect -419 -731 -385 -705
rect 1177 -731 1211 -705
rect -419 -765 -359 -731
rect 1151 -765 1211 -731
<< psubdiffcont >>
rect -359 695 1151 729
rect -419 -705 -385 669
rect 1177 -705 1211 669
rect -359 -765 1151 -731
<< poly >>
rect 217 525 482 560
rect 58 -74 657 0
rect 217 -632 486 -599
<< locali >>
rect -419 695 -359 729
rect 1151 695 1211 729
rect -419 669 -385 695
rect -419 -731 -385 -705
rect 1177 669 1211 695
rect 1177 -731 1211 -705
rect -419 -765 -359 -731
rect 1151 -765 1211 -731
<< viali >>
rect 272 729 306 730
rect 272 695 306 729
rect 272 694 306 695
rect 404 -731 448 -730
rect 404 -765 448 -731
rect 404 -766 448 -765
<< metal1 >>
rect 266 730 312 742
rect 266 694 272 730
rect 306 694 312 730
rect 266 682 312 694
rect -234 487 -198 561
rect -237 84 55 486
rect 272 458 306 682
rect 877 488 908 566
rect 659 476 915 488
rect -236 83 52 84
rect 6 56 52 83
rect 6 10 116 56
rect 270 -30 304 120
rect 394 100 404 476
rect 456 100 466 476
rect 651 100 661 476
rect 713 100 915 476
rect 659 89 915 100
rect 270 -32 424 -30
rect 270 -66 446 -32
rect -198 -172 53 -161
rect -198 -548 2 -172
rect 54 -548 64 -172
rect -198 -561 53 -548
rect 251 -549 261 -173
rect 313 -549 323 -173
rect 410 -200 446 -66
rect 619 -123 707 -88
rect 666 -160 707 -123
rect -193 -639 -160 -561
rect 410 -724 444 -534
rect 663 -560 912 -160
rect 871 -592 906 -560
rect 870 -638 906 -592
rect 392 -730 460 -724
rect 392 -766 404 -730
rect 448 -766 460 -730
rect 392 -772 460 -766
<< via1 >>
rect 404 100 456 476
rect 661 100 713 476
rect 2 -548 54 -172
rect 261 -549 313 -173
<< metal2 >>
rect 404 476 456 486
rect 400 100 404 146
rect 400 94 456 100
rect 659 476 715 486
rect 400 -30 450 94
rect 659 90 715 100
rect 260 -66 450 -30
rect 0 -172 56 -162
rect 260 -173 320 -66
rect 260 -176 261 -173
rect 0 -558 56 -548
rect 313 -176 320 -173
rect 261 -559 313 -549
<< via2 >>
rect 659 100 661 476
rect 661 100 713 476
rect 713 100 715 476
rect 0 -548 2 -172
rect 2 -548 54 -172
rect 54 -548 56 -172
<< metal3 >>
rect 649 476 725 481
rect 649 100 659 476
rect 715 100 725 476
rect 649 95 725 100
rect 658 -8 725 95
rect -9 -75 725 -8
rect -9 -167 58 -75
rect -10 -172 66 -167
rect -10 -548 0 -172
rect 56 -548 66 -172
rect -10 -553 66 -548
use sky130_fd_pr__nfet_01v8_7CP4KT  sky130_fd_pr__nfet_01v8_7CP4KT_0
timestamp 1729233293
transform 1 0 849 0 1 319
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_46AAJJ  sky130_fd_pr__nfet_01v8_46AAJJ_0
timestamp 1729224535
transform 1 0 158 0 1 288
box -158 -288 158 288
use sky130_fd_pr__nfet_01v8_46AAJJ  sky130_fd_pr__nfet_01v8_46AAJJ_1
timestamp 1729224535
transform 1 0 158 0 1 -360
box -158 -288 158 288
use sky130_fd_pr__nfet_01v8_46AAJJ  sky130_fd_pr__nfet_01v8_46AAJJ_2
timestamp 1729224535
transform 1 0 557 0 1 288
box -158 -288 158 288
use sky130_fd_pr__nfet_01v8_46AAJJ  sky130_fd_pr__nfet_01v8_46AAJJ_3
timestamp 1729224535
transform 1 0 557 0 1 -361
box -158 -288 158 288
use sky130_fd_pr__nfet_01v8_L2VWCK  sky130_fd_pr__nfet_01v8_L2VWCK_0
timestamp 1729233293
transform 1 0 -132 0 1 -392
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_LG94FM  sky130_fd_pr__nfet_01v8_LG94FM_0
timestamp 1729233293
transform 1 0 -170 0 1 318
box -73 -257 73 257
use sky130_fd_pr__nfet_01v8_SCJFGL  sky130_fd_pr__nfet_01v8_SCJFGL_0
timestamp 1729233293
transform 1 0 867 0 1 -387
box -73 -257 73 257
<< labels >>
flabel metal1 30 54 30 54 0 FreeSans 1600 0 0 0 D3
port 0 nsew
flabel metal2 422 24 422 24 0 FreeSans 1600 0 0 0 RS
port 1 nsew
flabel metal3 692 34 692 34 0 FreeSans 1600 0 0 0 D4
port 2 nsew
flabel metal1 288 604 288 604 0 FreeSans 1600 0 0 0 GND
port 3 nsew
<< end >>
