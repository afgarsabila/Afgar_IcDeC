magic
tech sky130A
magscale 1 2
timestamp 1729067780
<< viali >>
rect -3 -1158 1050 -1088
rect 12 -2231 1050 -2149
<< metal1 >>
rect -18 -1088 1072 -1038
rect -18 -1158 -3 -1088
rect 1050 -1158 1072 -1088
rect -18 -1160 1072 -1158
rect -15 -1164 1062 -1160
rect 166 -1679 176 -1627
rect 228 -1679 238 -1627
rect 314 -1672 510 -1637
rect 630 -1672 826 -1637
rect 892 -1677 902 -1625
rect 954 -1677 964 -1625
rect 0 -2143 1054 -2139
rect 0 -2149 1062 -2143
rect 0 -2231 12 -2149
rect 1050 -2231 1062 -2149
rect 0 -2237 1062 -2231
rect 0 -2241 1054 -2237
<< via1 >>
rect 176 -1679 228 -1627
rect 902 -1677 954 -1625
<< metal2 >>
rect 176 -1625 228 -1617
rect 166 -1627 228 -1625
rect 902 -1625 954 -1615
rect 166 -1677 176 -1627
rect 228 -1677 902 -1627
rect 954 -1677 964 -1625
rect 228 -1679 954 -1677
rect 176 -1689 228 -1679
rect 902 -1687 954 -1679
use inverterspice  x1
timestamp 1729049045
transform 1 0 -1146 0 1 -2585
box 1146 373 1568 1499
use inverterspice  x2
timestamp 1729049045
transform 1 0 -830 0 1 -2585
box 1146 373 1568 1499
use inverterspice  x3
timestamp 1729049045
transform 1 0 -514 0 1 -2585
box 1146 373 1568 1499
<< labels >>
flabel viali 39 -1139 39 -1139 0 FreeSans 320 0 0 0 vdd
port 0 nsew
flabel viali 309 -2222 309 -2222 0 FreeSans 320 0 0 0 gnd
port 1 nsew
flabel via1 930 -1653 930 -1653 0 FreeSans 320 0 0 0 out
port 2 nsew
<< end >>
